-- PLL_Reconfig.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PLL_Reconfig is
	port (
		mgmt_clk          : in  std_logic                     := '0';             --          mgmt_clk.clk
		mgmt_reset        : in  std_logic                     := '0';             --        mgmt_reset.reset
		mgmt_waitrequest  : out std_logic;                                        -- mgmt_avalon_slave.waitrequest
		mgmt_read         : in  std_logic                     := '0';             --                  .read
		mgmt_write        : in  std_logic                     := '0';             --                  .write
		mgmt_readdata     : out std_logic_vector(31 downto 0);                    --                  .readdata
		mgmt_address      : in  std_logic_vector(5 downto 0)  := (others => '0'); --                  .address
		mgmt_writedata    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .writedata
		reconfig_to_pll   : out std_logic_vector(63 downto 0);                    --   reconfig_to_pll.reconfig_to_pll
		reconfig_from_pll : in  std_logic_vector(63 downto 0) := (others => '0')  -- reconfig_from_pll.reconfig_from_pll
	);
end entity PLL_Reconfig;

architecture rtl of PLL_Reconfig is
	component altera_pll_reconfig_top is
		generic (
			device_family       : string  := "";
			ENABLE_MIF          : boolean := false;
			MIF_FILE_NAME       : string  := "";
			ENABLE_BYTEENABLE   : boolean := false;
			BYTEENABLE_WIDTH    : integer := 4;
			RECONFIG_ADDR_WIDTH : integer := 6;
			RECONFIG_DATA_WIDTH : integer := 32;
			reconf_width        : integer := 64;
			WAIT_FOR_LOCK       : boolean := true
		);
		port (
			mgmt_clk          : in  std_logic                     := 'X';             -- clk
			mgmt_reset        : in  std_logic                     := 'X';             -- reset
			mgmt_waitrequest  : out std_logic;                                        -- waitrequest
			mgmt_read         : in  std_logic                     := 'X';             -- read
			mgmt_write        : in  std_logic                     := 'X';             -- write
			mgmt_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			mgmt_address      : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			mgmt_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reconfig_to_pll   : out std_logic_vector(63 downto 0);                    -- reconfig_to_pll
			reconfig_from_pll : in  std_logic_vector(63 downto 0) := (others => 'X'); -- reconfig_from_pll
			mgmt_byteenable   : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- byteenable
		);
	end component altera_pll_reconfig_top;

begin

	pll_reconfig_inst : component altera_pll_reconfig_top
		generic map (
			device_family       => "Cyclone V",
			ENABLE_MIF          => false,
			MIF_FILE_NAME       => "",
			ENABLE_BYTEENABLE   => false,
			BYTEENABLE_WIDTH    => 4,
			RECONFIG_ADDR_WIDTH => 6,
			RECONFIG_DATA_WIDTH => 32,
			reconf_width        => 64,
			WAIT_FOR_LOCK       => true
		)
		port map (
			mgmt_clk          => mgmt_clk,          --          mgmt_clk.clk
			mgmt_reset        => mgmt_reset,        --        mgmt_reset.reset
			mgmt_waitrequest  => mgmt_waitrequest,  -- mgmt_avalon_slave.waitrequest
			mgmt_read         => mgmt_read,         --                  .read
			mgmt_write        => mgmt_write,        --                  .write
			mgmt_readdata     => mgmt_readdata,     --                  .readdata
			mgmt_address      => mgmt_address,      --                  .address
			mgmt_writedata    => mgmt_writedata,    --                  .writedata
			reconfig_to_pll   => reconfig_to_pll,   --   reconfig_to_pll.reconfig_to_pll
			reconfig_from_pll => reconfig_from_pll, -- reconfig_from_pll.reconfig_from_pll
			mgmt_byteenable   => "0000"             --       (terminated)
		);

end architecture rtl; -- of PLL_Reconfig
